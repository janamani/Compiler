module SARFastVerilog(Clock, Reset, Inc, Dcr, Compare, DataOut,
     ClockCmp, StateP, SAROut);
  input Clock, Reset, Inc, Dcr, Compare;
  input [7:0] DataOut;
  output ClockCmp;
  output [1:0] StateP;
  output [7:0] SAROut;
  wire Clock, Reset, Inc, Dcr, Compare;
  wire [7:0] DataOut;
  wire ClockCmp;
  wire [1:0] StateP;
  wire [7:0] SAROut;
  wire [7:0] SAR;
  wire [7:0] TempSAR;
  wire [1:0] CheckID;
  wire N0, N1, N3, N4, N6, N7, N8, N9;
  wire N10, N11, N12, N13, N14, N15, N17, N18;
  wire N19, N20, N21, N22, N23, N24, N25, N26;
  wire N27, N28, N29, N30, N31, N32, N33, N35;
  wire N36, N37, N38, N39, N40, N42, N43, N44;
  wire N45, N46, N47, N48, N49, N50, N51, N52;
  wire N53, N54, N55, N56, N57, N58, N59, N60;
  wire N61, N62, N63, N64, N65, N66, N67, N68;
  wire N69, N70, N71, N72, N73, N74, N75, N76;
  wire N77, N79, N80, N81, N82, N83, N84, N85;
  wire N86, N87, N88, N89, N90, N91, N92, N93;
  wire N94, N95, N96, N97, N98, N99, N100, N101;
  wire N102, N103, N104, N105, N106, N107, N108, N109;
  wire N110, N111, N112, N118, N119, N120, N121, N122;
  wire N123, N134, N135, N137, N138, N139, N140, N141;
  wire N142, N143, N144, N145, N146, N147, N149, N150;
  wire N159, N160, N161;
  INV1S g2485(.I (N150), .O (N112));
  INV1S g2486(.I (N123), .O (N135));
  OR2 g2483(.I1 (StateP[0]), .I2 (StateP[1]), .O (N123));
  NR2 g3022(.I1 (Reset), .I2 (N111), .O (SAROut[0]));
  INV1S g3023(.I (N111), .O (N144));
  NR2 g3024(.I1 (SAR[0]), .I2 (TempSAR[0]), .O (N111));
  QDFFRBS \SAR_reg[0] (.RB (N4), .CK (Clock), .D (N110), .Q (SAR[0]));
  AO222 g3026(.A1 (N85), .A2 (SAR[1]), .B1 (N98), .B2 (N86), .C1 (N87), .C2 (N101), .O (N110));
  AN2 g3027(.I1 (N143), .I2 (N4), .O (SAROut[1]));
  OR2 g3028(.I1 (SAR[1]), .I2 (TempSAR[1]), .O (N143));
  QDFFRBS \SAR_reg[1] (.RB (N4), .CK (Clock), .D (N109), .Q (SAR[1]));
  AO222 g3030(.A1 (N85), .A2 (SAR[2]), .B1 (N98), .B2 (N77), .C1 (N87), .C2 (N100), .O (N109));
  AN2 g3031(.I1 (N142), .I2 (N4), .O (SAROut[2]));
  OR2 g3032(.I1 (SAR[2]), .I2 (TempSAR[2]), .O (N142));
  QDFFRBS \SAR_reg[2] (.RB (N4), .CK (Clock), .D (N108), .Q (SAR[2]));
  AO222 g3034(.A1 (N85), .A2 (SAR[3]), .B1 (N98), .B2 (DataOut[2]), .C1 (N87), .C2 (N99), .O (N108));
  AN2 g3035(.I1 (N141), .I2 (N4), .O (SAROut[3]));
  OR2 g3036(.I1 (SAR[3]), .I2 (TempSAR[3]), .O (N141));
  QDFFRBS \SAR_reg[3] (.RB (N4), .CK (Clock), .D (N107), .Q (SAR[3]));
  ND2 g3038(.I1 (N106), .I2 (N97), .O (N107));
  AN2 g3039(.I1 (N140), .I2 (N4), .O (SAROut[4]));
  AOI22S g3040(.A1 (N85), .A2 (SAR[4]), .B1 (N87), .B2 (N96), .O (N106));
  OR2 g3041(.I1 (SAR[4]), .I2 (TempSAR[4]), .O (N140));
  QDFFRBS \SAR_reg[4] (.RB (N4), .CK (Clock), .D (N105), .Q (SAR[4]));
  AO222 g3043(.A1 (N85), .A2 (SAR[5]), .B1 (N94), .B2 (DataOut[4]), .C1 (N87), .C2 (N92), .O (N105));
  AN2 g3044(.I1 (N139), .I2 (N4), .O (SAROut[5]));
  OR2 g3045(.I1 (SAR[5]), .I2 (TempSAR[5]), .O (N139));
  QDFFRBS \SAR_reg[5] (.RB (N4), .CK (Clock), .D (N104), .Q (SAR[5]));
  ND2 g3047(.I1 (N103), .I2 (N93), .O (N104));
  AN2 g3048(.I1 (N138), .I2 (N4), .O (SAROut[6]));
  AOI22S g3049(.A1 (N85), .A2 (SAR[6]), .B1 (N87), .B2 (N88), .O (N103));
  OR2 g3050(.I1 (SAR[6]), .I2 (TempSAR[6]), .O (N138));
  QDFFRBS \SAR_reg[6] (.RB (N4), .CK (Clock), .D (N102), .Q (SAR[6]));
  AO222 g3052(.A1 (N85), .A2 (SAR[7]), .B1 (N90), .B2 (DataOut[6]), .C1 (N87), .C2 (N84), .O (N102));
  AN2 g3053(.I1 (N137), .I2 (N4), .O (SAROut[7]));
  INV1S g3054(.I (N101), .O (N147));
  NR2 g3055(.I1 (DataOut[0]), .I2 (N150), .O (N101));
  OR2 g3056(.I1 (SAR[7]), .I2 (TempSAR[7]), .O (N137));
  NR2 g3057(.I1 (DataOut[1]), .I2 (N119), .O (N100));
  OR2B1S g3058(.I1 (N119), .B1 (DataOut[1]), .O (N150));
  QDFFRBS \SAR_reg[7] (.RB (N4), .CK (Clock), .D (N95), .Q (SAR[7]));
  NR2 g3060(.I1 (DataOut[2]), .I2 (N120), .O (N99));
  OR2B1S g3061(.I1 (N120), .B1 (DataOut[2]), .O (N119));
  AN3B2S g3062(.I1 (N94), .B1 (DataOut[4]), .B2 (DataOut[3]), .O (N98));
  ND3 g3063(.I1 (N94), .I2 (N81), .I3 (DataOut[3]), .O (N97));
  NR2 g3064(.I1 (DataOut[3]), .I2 (N121), .O (N96));
  ND2 g3065(.I1 (N91), .I2 (DataOut[3]), .O (N120));
  NR2 g3066(.I1 (N134), .I2 (N89), .O (N95));
  AN3B2S g3067(.I1 (N90), .B1 (DataOut[6]), .B2 (DataOut[5]), .O (N94));
  ND3 g3068(.I1 (N90), .I2 (N82), .I3 (DataOut[5]), .O (N93));
  NR2 g3069(.I1 (DataOut[4]), .I2 (N122), .O (N92));
  INV1S g3070(.I (N91), .O (N121));
  NR2 g3071(.I1 (N81), .I2 (N122), .O (N91));
  NR3 g3072(.I1 (DataOut[7]), .I2 (N146), .I3 (N134), .O (N90));
  MUX2 g3073(.S (DataOut[7]), .A (N145), .B (N146), .O (N89));
  ND2 g3074(.I1 (N118), .I2 (DataOut[5]), .O (N122));
  NR2 g3075(.I1 (DataOut[5]), .I2 (N83), .O (N88));
  NR2 g3076(.I1 (N145), .I2 (N134), .O (N87));
  NR3 g3077(.I1 (Clock), .I2 (N135), .I3 (Reset), .O (ClockCmp));
  AN3B2S g3078(.I1 (DataOut[0]), .B1 (DataOut[2]), .B2 (DataOut[1]), .O (N86));
  AN2 g3079(.I1 (N79), .I2 (StateP[1]), .O (N85));
  ND2 g3080(.I1 (N80), .I2 (CheckID[0]), .O (N146));
  OR2 g3081(.I1 (CheckID[0]), .I2 (N80), .O (N145));
  OR2 g3082(.I1 (StateP[1]), .I2 (N79), .O (N134));
  AN2 g3083(.I1 (N82), .I2 (DataOut[7]), .O (N84));
  INV1S g3084(.I (N83), .O (N118));
  ND2S g3085(.I1 (DataOut[6]), .I2 (DataOut[7]), .O (N83));
  ND2 g3087(.I1 (DataOut[1]), .I2 (DataOut[6]), .O (N149));
  INV1S g3088(.I (DataOut[6]), .O (N82));
  INV1S g3089(.I (DataOut[4]), .O (N81));
  INV1S g3093(.I (Reset), .O (N4));
  AN2B1S g2(.I1 (DataOut[1]), .B1 (DataOut[2]), .O (N77));
  DFFRBN \TempSAR_reg[0] (.RB (N4), .CK (Clock), .D (N66), .Q (TempSAR[0]), .QB (N160));
  QDFFRBN \TempSAR_reg[1] (.RB (N4), .CK (Clock), .D (N74), .Q (TempSAR[1]));
  QDFFRBN \TempSAR_reg[6] (.RB (N4), .CK (Clock), .D (N73), .Q (TempSAR[6]));
  QDFFRBN \TempSAR_reg[3] (.RB (N4), .CK (Clock), .D (N72), .Q (TempSAR[3]));
  QDFFRBN \TempSAR_reg[2] (.RB (N4), .CK (Clock), .D (N75), .Q (TempSAR[2]));
  QDFFRBN \TempSAR_reg[4] (.RB (N4), .CK (Clock), .D (N71), .Q (TempSAR[4]));
  QDFFRBN \TempSAR_reg[5] (.RB (N4), .CK (Clock), .D (N76), .Q (TempSAR[5]));
  QDFFRBN \TempSAR_reg[7] (.RB (N4), .CK (Clock), .D (N70), .Q (TempSAR[7]));
  DFFSBN \StateP_reg[0] (.SB (N4), .CK (Clock), .D (N69), .Q (StateP[0]), .QB (N79));
  ND2 g3624(.I1 (N68), .I2 (N26), .O (N76));
  ND3 g3625(.I1 (N57), .I2 (N64), .I3 (N27), .O (N75));
  AO12 g3626(.A1 (N67), .B1 (N8), .B2 (N143), .O (N74));
  AO222 g3627(.A1 (N8), .A2 (N138), .B1 (N60), .B2 (TempSAR[6]), .C1 (N36), .C2 (N161), .O (N73));
  AO222 g3628(.A1 (N8), .A2 (N141), .B1 (N62), .B2 (TempSAR[3]), .C1 (N19), .C2 (N55), .O (N72));
  AO222 g3629(.A1 (N8), .A2 (N140), .B1 (N62), .B2 (TempSAR[4]), .C1 (N19), .C2 (N54), .O (N71));
  ND3 g3630(.I1 (N65), .I2 (N50), .I3 (N25), .O (N70));
  OAI12S g3631(.A1 (N4), .B1 (N61), .B2 (N56), .O (N69));
  AOI112S g3632(.A1 (N53), .B1 (N40), .C1 (N62), .C2 (TempSAR[5]), .O (N68));
  MOAI1S g3633(.A1 (N20), .A2 (N147), .B1 (N62), .B2 (TempSAR[1]), .O (N67));
  MOAI1S g3634(.A1 (N59), .A2 (N160), .B1 (N8), .B2 (N144), .O (N66));
  OAI12S g3635(.A1 (TempSAR[7]), .B1 (N58), .B2 (N0), .O (N65));
  OA13S g3636(.A1 (N63), .B1 (N20), .B2 (N43), .B3 (N119), .O (N64));
  ND2 g3637(.I1 (N58), .I2 (TempSAR[2]), .O (N63));
  AO12 g3638(.A1 (N58), .B1 (N7), .B2 (N42), .O (N62));
  AOI112S g3639(.A1 (N52), .B1 (N134), .C1 (N146), .C2 (N42), .O (N61));
  AO12 g3640(.A1 (N58), .B1 (N7), .B2 (N118), .O (N60));
  AOI13HS g3641(.A1 (N58), .B1 (N7), .B2 (N112), .B3 (DataOut[0]), .O (N59));
  QDFFRBN \CheckID_reg[0] (.RB (N4), .CK (Clock), .D (N49), .Q (CheckID[0]));
  DFFSBN \StateP_reg[1] (.SB (N4), .CK (Clock), .D (N51), .Q (StateP[1]), .QB (N3));
  ND2 g3645(.I1 (N45), .I2 (N46), .O (N58));
  ND3 g3646(.I1 (N48), .I2 (N43), .I3 (DataOut[2]), .O (N57));
  OAI112S g3647(.A1 (N21), .B1 (N11), .C1 (N3), .C2 (N31), .O (N56));
  MOAI1S g3648(.A1 (N120), .A2 (N159), .B1 (N43), .B2 (N38), .O (N55));
  OAI22S g3649(.A1 (N122), .A2 (N44), .B1 (N121), .B2 (N15), .O (N54));
  AOI112S g3650(.A1 (N35), .B1 (N14), .C1 (N33), .C2 (DataOut[4]), .O (N53));
  OA12 g3651(.A1 (N145), .B1 (N146), .B2 (N30), .O (N52));
  AO12 g3652(.A1 (Reset), .B1 (N123), .B2 (N11), .O (N51));
  OAI112S g3653(.A1 (N19), .B1 (DataOut[7]), .C1 (N39), .C2 (N28), .O (N50));
  AO22 g3654(.A1 (N18), .A2 (CheckID[0]), .B1 (N6), .B2 (Dcr), .O (N49));
  OAI22S g3655(.A1 (N120), .A2 (N37), .B1 (N24), .B2 (N149), .O (N48));
  AO22 g3656(.A1 (N18), .A2 (CheckID[1]), .B1 (N6), .B2 (Inc), .O (N47));
  OAI112S g3657(.A1 (N3), .B1 (CheckID[0]), .C1 (CheckID[1]), .C2 (N30), .O (N46));
  AOI112S g3658(.A1 (N6), .B1 (N17), .C1 (N7), .C2 (N80), .O (N45));
  OR2 g3659(.I1 (N29), .I2 (N33), .O (N44));
  NR2 g3660(.I1 (N1), .I2 (N39), .O (N43));
  NR2 g3661(.I1 (N29), .I2 (N32), .O (N42));
  NR3 g3663(.I1 (DataOut[0]), .I2 (N122), .I3 (N20), .O (N40));
  OR2B1S g3664(.I1 (N29), .B1 (DataOut[3]), .O (N39));
  AN2B1S g3665(.I1 (N28), .B1 (N121), .O (N38));
  ND2S g3666(.I1 (N19), .I2 (N149), .O (N37));
  INV1S g3667(.I (N35), .O (N36));
  ND2S g3668(.I1 (N19), .I2 (N118), .O (N35));
  INV1S g3670(.I (N32), .O (N33));
  OR3B2 g3671(.I1 (N28), .B1 (DataOut[7]), .B2 (DataOut[3]), .O (N32));
  AN4B1S g3672(.I1 (N23), .I2 (N13), .I3 (SAR[0]), .B1 (SAR[7]), .O (N31));
  AN4B1S g3673(.I1 (N22), .I2 (N10), .I3 (N1), .B1 (DataOut[0]), .O (N30));
  ND2 g3674(.I1 (N15), .I2 (DataOut[4]), .O (N29));
  ND3 g3675(.I1 (DataOut[1]), .I2 (DataOut[2]), .I3 (DataOut[6]), .O (N28));
  ND2 g3676(.I1 (N8), .I2 (N142), .O (N27));
  ND2 g3677(.I1 (N8), .I2 (N139), .O (N26));
  ND2 g3678(.I1 (N8), .I2 (N137), .O (N25));
  ND2S g3679(.I1 (N7), .I2 (TempSAR[2]), .O (N24));
  AN3B2S g3681(.I1 (N12), .B1 (SAR[1]), .B2 (SAR[2]), .O (N23));
  AN3B2S g3682(.I1 (N9), .B1 (DataOut[3]), .B2 (DataOut[6]), .O (N22));
  OR3 g3683(.I1 (Dcr), .I2 (Inc), .I3 (N123), .O (N21));
  INV1S g3684(.I (N20), .O (N19));
  ND3 g3685(.I1 (N7), .I2 (StateP[0]), .I3 (CheckID[1]), .O (N20));
  MOAI1S g3686(.A1 (N3), .A2 (StateP[0]), .B1 (N3), .B2 (StateP[0]), .O (N18));
  NR2 g3687(.I1 (Compare), .I2 (N3), .O (N17));
  INV1S g3689(.I (N14), .O (N15));
  ND2S g3690(.I1 (DataOut[5]), .I2 (DataOut[0]), .O (N14));
  NR2 g3691(.I1 (SAR[6]), .I2 (SAR[5]), .O (N13));
  NR2 g3692(.I1 (SAR[4]), .I2 (SAR[3]), .O (N12));
  ND2 g3693(.I1 (StateP[0]), .I2 (StateP[1]), .O (N11));
  NR2 g3694(.I1 (DataOut[4]), .I2 (DataOut[2]), .O (N10));
  NR2 g3695(.I1 (DataOut[1]), .I2 (DataOut[5]), .O (N9));
  AN2 g3696(.I1 (StateP[1]), .I2 (Compare), .O (N8));
  NR2 g3698(.I1 (CheckID[0]), .I2 (StateP[1]), .O (N7));
  NR2 g3699(.I1 (StateP[1]), .I2 (StateP[0]), .O (N6));
  INV1S g3723(.I (DataOut[7]), .O (N1));
  AN2B1S g3094(.I1 (N7), .B1 (N1), .O (N0));
  INV1S g3725(.I (N29), .O (N159));
  DFFRBN \CheckID_reg[1] (.RB (N4), .CK (Clock), .D (N47), .Q (CheckID[1]), .QB (N80));


  OR3B2 g3730(.I1 (N39), .B1 (DataOut[2]), .B2 (DataOut[1]), .O (N161));
endmodule

